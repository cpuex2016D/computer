parameter INST_WIDTH = 32;
parameter REG_WIDTH = 5;
parameter ROB_WIDTH = 4;
