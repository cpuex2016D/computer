`include "common.vh"

module add_sub_tb;
	logic clk = 0;
	unit_if i();
	add_sub add_sub(.*);
	localparam OP_ADD     = 6'b000000;
	localparam OP_ADDI    = 6'b000001;
	localparam OP_SUB     = 6'b000010;
	localparam OP_SUBI    = 6'b000011;
	localparam OP_SL2ADD  = 6'b000100;
	localparam OP_SL2ADDI = 6'b000101;

	always #(0.5) clk <= !clk;

	initial begin
		i.inst.bits <= {OP_ADD, 5'd0, 5'd0, 5'd0, 11'd0};
		i.read[0].valid <= 1;
		i.read[0].tag <= {ROB_WIDTH{1'bx}};
		i.read[0].data <= 2;
		i.read[1].valid <= 1;
		i.read[1].tag <= {ROB_WIDTH{1'bx}};
		i.read[1].data <= 3;
		i.new_tag <= 8;
		i.cdb.valid <= 0;
		i.cdb.tag <= {ROB_WIDTH{1'bx}};
		i.cdb.data <= 32'bx;
		i.req.ready <= 1;
		#1;
		i.inst.bits <= {OP_ADDI, 5'd0, 5'd0, 16'd1};
		i.read[0].valid <= 0;
		i.read[0].tag <= 0;
		i.read[0].data <= 32'bx;
		i.read[1].valid <= 1'bx;
		i.read[1].tag <= {ROB_WIDTH{1'bx}};
		i.read[1].data <= 32'bx;
		i.new_tag <= 9;
		i.cdb.valid <= 0;
		i.cdb.tag <= {ROB_WIDTH{1'bx}};
		i.cdb.data <= 32'bx;
		i.req.ready <= 1;
		#1;
		i.inst.bits <= 32'hffffffff;
		i.read[0].valid <= 1'bx;
		i.read[0].tag <= {ROB_WIDTH{1'bx}};
		i.read[0].data <= 32'bx;
		i.read[1].valid <= 1'bx;
		i.read[1].tag <= {ROB_WIDTH{1'bx}};
		i.read[1].data <= 32'bx;
		i.new_tag <= 10;
		i.cdb.valid <= 1;
		i.cdb.tag <= 0;
		i.cdb.data <= 10;
		i.req.ready <= 1;
		#1;
		i.inst.bits <= {OP_SL2ADDI, 5'd0, 5'd0, 16'd1};
		i.read[0].valid <= 1;
		i.read[0].tag <= {ROB_WIDTH{1'bx}};
		i.read[0].data <= 1;
		i.read[1].valid <= 1'bx;
		i.read[1].tag <= {ROB_WIDTH{1'bx}};
		i.read[1].data <= 32'bx;
		i.new_tag <= 11;
		i.cdb.valid <= 0;
		i.cdb.tag <= {ROB_WIDTH{1'bx}};
		i.cdb.data <= 32'bx;
		i.req.ready <= 1;

		#1;
		i.inst.bits <= {OP_ADD, 5'd0, 5'd0, 5'd0, 11'd0};
		i.read[0].valid <= 1;
		i.read[0].tag <= {ROB_WIDTH{1'bx}};
		i.read[0].data <= 2;
		i.read[1].valid <= 1;
		i.read[1].tag <= {ROB_WIDTH{1'bx}};
		i.read[1].data <= 3;
		i.new_tag <= 12;
		i.cdb.valid <= 0;
		i.cdb.tag <= {ROB_WIDTH{1'bx}};
		i.cdb.data <= 32'bx;
		i.req.ready <= 0;
		#1;
		i.inst.bits <= {OP_ADDI, 5'd0, 5'd0, 16'd1};
		i.read[0].valid <= 0;
		i.read[0].tag <= 0;
		i.read[0].data <= 32'bx;
		i.read[1].valid <= 1'bx;
		i.read[1].tag <= {ROB_WIDTH{1'bx}};
		i.read[1].data <= 32'bx;
		i.new_tag <= 13;
		i.cdb.valid <= 0;
		i.cdb.tag <= {ROB_WIDTH{1'bx}};
		i.cdb.data <= 32'bx;
		i.req.ready <= 0;
		#1;
		i.inst.bits <= 32'hffffffff;
		i.read[0].valid <= 1'bx;
		i.read[0].tag <= {ROB_WIDTH{1'bx}};
		i.read[0].data <= 32'bx;
		i.read[1].valid <= 1'bx;
		i.read[1].tag <= {ROB_WIDTH{1'bx}};
		i.read[1].data <= 32'bx;
		i.new_tag <= 14;
		i.cdb.valid <= 1;
		i.cdb.tag <= 0;
		i.cdb.data <= 10;
		i.req.ready <= 0;
		#1;
		i.inst.bits <= {OP_SL2ADDI, 5'd0, 5'd0, 16'd1};
		i.read[0].valid <= 1;
		i.read[0].tag <= {ROB_WIDTH{1'bx}};
		i.read[0].data <= 1;
		i.read[1].valid <= 1'bx;
		i.read[1].tag <= {ROB_WIDTH{1'bx}};
		i.read[1].data <= 32'bx;
		i.new_tag <= 15;
		i.cdb.valid <= 0;
		i.cdb.tag <= {ROB_WIDTH{1'bx}};
		i.cdb.data <= 32'bx;
		i.req.ready <= 0;
	end
endmodule
