import my_package::*;
